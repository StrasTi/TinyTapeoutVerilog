module n_bit_alu(
    input a_i,
    input b_i,
    input [3:0] f_i,
    output result_o,
    output carry_bit_o
);

endmodule
